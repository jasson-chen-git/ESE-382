---------------------------------------------------------------------------
----
--
-- Title : Design Task 5
-- Design : Sine Lookup Table
-- Author : Jason Chen
-- Company : 112515450
--
---------------------------------------------------------------------------
----
--
-- Description : Write a behavioral description for the sine table.
--
---------------------------------------------------------------------------
----
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;	

entity sine_table is
	port(
		addr : in std_logic_vector(6 downto 0);
		sine_val : out std_logic_vector(6 downto 0)
		);
end entity;

architecture behavioral of sine_table is
	type table_lookup is array (0 to 127) of std_logic_vector(6 downto 0);
	constant st : table_lookup := (
		"0000000", "0000001", "0000011", "0000100", "0000110", "0000111", 
		"0001001", "0001010", "0001100", "0001110", "0001111", "0010001", 
		"0010010", "0010100", "0010101", "0010111", "0011000", "0011010", 
		"0011100", "0011101", "0011111", "0100000", "0100010", "0100011", 
		"0100101", "0100110", "0101000", "0101001", "0101011", "0101100", 
		"0101110", "0101111", "0110000", "0110010", "0110011", "0110101", 
		"0110110", "0111000", "0111001", "0111010", "0111100", "0111101", 
		"0111111", "1000000", "1000001", "1000011", "1000100", "1000101", 
		"1000111", "1001000", "1001001", "1001010", "1001100", "1001101", 
		"1001110", "1001111", "1010001", "1010010", "1010011", "1010100", 
		"1010101", "1010111", "1011000", "1011001", "1011010", "1011011", 
		"1011100", "1011101", "1011110", "1011111", "1100000", "1100001", 
		"1100010", "1100011", "1100100", "1100101", "1100110", "1100111", 
		"1101000", "1101001", "1101010", "1101011", "1101100", "1101100", 
		"1101101", "1101110", "1101111", "1110000", "1110000", "1110001", 
		"1110010", "1110011", "1110011", "1110100", "1110101", "1110101", 
		"1110110", "1110110", "1110111", "1110111", "1111000", "1111001", 
		"1111001", "1111010", "1111010", "1111010", "1111011", "1111011", 
		"1111100", "1111100", "1111100", "1111101", "1111101", "1111101", 
		"1111110", "1111110", "1111110", "1111110", "1111111", "1111111", 
		"1111111", "1111111", "1111111", "1111111", "1111111", "1111111", 
		"1111111", "1111111"
		);
	begin		
		sine_val <= st(to_integer(unsigned(addr)));
end architecture;